package rst_agent_pkg;

	import uvm_pkg::*;

	typedef class agent_rst;
	typedef class config_rst;
	typedef class driver_rst;
	typedef class mon_rst;
	typedef class seq_item_rst;
	typedef class sequ_rst;
	typedef class sequencer_rst;

	`include "agent_rst.sv"
	`include "config_rst.sv"
	`include "driver_rst.sv"
	`include "mon_rst.sv"
	`include "seq_item_rst.sv"
	`include "sequ_rst.sv"
	`include "sequencer_rst.sv"

endpackage