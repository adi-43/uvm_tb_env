`ifndef INTF_RST
    `define INTF_RST

interface intf_rst();
    
    bit rst_in;
    bit rst_out;

endinterface

`endif
